%!PS-Adobe-3.0 EPSF-3.0
%%Title: ha2.ckt
%%Creator: XCircuit v3.6 rev78
%%CreationDate: Sat Dec 15 15:02:30 2007
%%Pages: 1
%%BoundingBox: 68 68 652 354
%%DocumentNeededResources: font Helvetica Times-Roman Symbol 
%%EndComments
%%BeginProlog
%
%  PostScript prolog for output from xcircuit
%  Version: 3.3
%
%  Electrical circuit (and otherwise general) drawing program
%
%  Written by Tim Edwards 8/5/93--7/13/05  (tim.edwards@multigig.com)
%  The Johns Hopkins University (1993-2004)
%  MultiGiG, Inc. (2004-present)
%
%%BeginResource: procset XCIRCproc 3.3 0
%
% supporting definitions --- these are the primary xcircuit types.

/XCIRCsave save def
/topmat matrix currentmatrix def

/fontslant { /slant exch def [1 0 slant 1 0 0] 
    exch findfont exch makefont dup length dict /ndict exch def
    { 1 index /FID ne { ndict 3 1 roll put } { pop pop } ifelse } forall
    ndict definefont pop} def
/ul { dup type /stringtype eq showflag 1 eq and { gsave 
   currentpoint topmat setmatrix 0 0 moveto 2 index stringwidth pop (_)
   false charpath flattenpath pathbbox grestore exch pop 1 index
   sub setlinewidth exch pop currentpoint 3 -1 roll add moveto 0
   rlineto stroke moveto } if } def
/ol { dup type /stringtype eq showflag 1 eq and { gsave gsave
   currentpoint topmat setmatrix 2 index stringwidth pop 3 index
   true charpath flattenpath pathbbox grestore exch pop
   exch pop topmat setmatrix (_) true charpath pathbbox grestore
   exch pop 1 index sub setlinewidth exch pop currentpoint
   exch 4 1 roll exch sub add moveto pop 0 rlineto stroke
   moveto } if } def
/stW { gsave currentpoint newpath moveto true charpath flattenpath
	pathbbox pop exch pop sub grestore } def
/Ts {mark Tabs aload pop counttomark 1 add array astore /Tabs exch def Tabs
	0 currentpoint pop put} def
/Tbn {mark Tabs aload pop counttomark dup 2 add 1 roll cleartomark 1 sub} def
/Tb { 0 1 Tbn {Tabs exch get dup currentpoint pop lt
	{currentpoint exch pop moveto exit} {pop} ifelse } for } def
/Tf { Tbn -1 0 {Tabs exch get dup currentpoint pop gt
	{currentpoint exch pop moveto exit} {pop} ifelse } for } def
/qS { (aa) stW (a a) stW sub 4 div 0 Kn } def
/hS { qS qS } def
/pspc 0 def
/cf0 { scalefont setfont } bind def
/Kn { dup kY add /kY exch def rmoveto } bind def
/ss { /fscale fscale 0.67 mul def currentfont 0.67 cf0 0 fscale0 fscale mul
	0.33 mul neg Kn} def
/Ss { /fscale fscale 0.67 mul def currentfont 0.67 cf0 0 fscale0 fscale mul
	0.67 mul Kn } def
/ns { 0 kY neg Kn /kY 0 def /fscale 1.0 def xfont0 1.0 cf0 } def
/CR { ns 0 /Bline Bline fscale0 neg add def Bline moveto } def
/cf { dup type /realtype ne {1.0} if exch findfont exch kY 0 eq
	{ 40 mul dup /fscale0 exch def cf0 /xfont0 currentfont def}
	{fscale0 mul fscale mul cf0} ifelse } def
/ctmk { counttomark dup 2 add -1 roll pop } bind def
/label { gsave translate 0 0 moveto dup scale neg /rotval exch def
	/just exch def just 384 and 0 gt {/mshow {pop} def} {/mshow {show}
	def} ifelse just 16 and 0 gt {gsave rotval rotate 0 1 dtransform
	gsave pagemat setmatrix idtransform exch grestore 1 0 dtransform
	gsave pagemat setmatrix idtransform exch grestore dup abs 1e-9 lt
	{pop mul 0 gt} {3 1 roll pop pop 0 lt} ifelse grestore {-1 /rotval
	rotval neg def /just just dup 3 and 1 ne {3 xor} if def} {1} ifelse
	exch -1e-9 lt {-1 /rotval rotval neg def /just just dup 12 and
	4 ne {12 xor} if def} {1} ifelse scale } if /showflag 0 def
	/fspc pspc def /Bline 0 def /Tabs 0 array def /fscale 1.0 def
	/kY 0 def gsave dup 1 add copy 0 exch 1 0 dtransform exch atan rotate
	{exch dup type /stringtype eq {true charpath flattenpath} {dup type
	/arraytype eq {exec} {12 string cvs true charpath flattenpath} ifelse}
	ifelse} repeat pop pathbbox grestore 3 -1 roll pop 3 1 roll just
	1 and 0 gt {just 2 and 0 gt {exch pop neg fspc sub} {exch sub 0.5
	mul neg} ifelse} {pop neg fspc add} ifelse exch Bline exch just 4
	and 0 gt {just 8 and 0 gt {exch pop neg fspc sub} {add 0.5 mul neg}
	ifelse} {pop neg fspc add} ifelse rotval rotate Kn currentpoint
	translate /showflag 1 def /Bline 0 def /Tabs 0 array def /fscale
	1.0 def /kY 0 def {dup type /stringtype eq {mshow} {dup type
	/arraytype eq {exec} {12 string cvs mshow} ifelse} ifelse} repeat
	grestore } def
/pinlabel { 4 index 32 and 0 ne hlevel 0 eq or { /pspc 10 def label
	/pspc 0 def } { pop pop pop pop pop {pop} repeat } ifelse } def
/pinglobal { pinlabel } def
/infolabel { pinlabel } def
/graphic { gsave 4 index cvx exec /DataSource get resetfile translate
	0 0 moveto neg rotate dup scale cvx exec image grestore } def

/scb { setrgbcolor } bind def  /sce { defColor aload pop scb } bind def
/cRedef {/defColor currentcolor 3 array astore def} def
/begingate {dup type /dicttype ne {1 dict} if begin	% default params
	dup type /dicttype ne {1 dict} if begin		% instanced params
	/hlevel hlevel 1 add def /defColor currentcolor sce 3 array
	astore def gsave sce translate 0 0 moveto neg rotate dup abs scale
	} bind def
/endgate { /hlevel hlevel 1 sub def grestore defColor aload pop cRedef
	scb end end} bind def

/hlevel 0 def
/tmpa [1 0 0 1 0 0] def
/gar {8 8 true tmpa {<c0 c0 00 00 0c 0c 00 00>} imagemask} bind
{8 8 true tmpa {<30 70 60 02 03 07 06 20>} imagemask} bind
{8 8 true tmpa {<0c 1e 1e 0c c0 e1 e1 c0>} imagemask} bind
{8 8 true tmpa {<0f 0f 0f 0f f0 f0 f0 f0>} imagemask} bind
{8 8 true tmpa {<3f f3 e1 e1 f3 3f 1e 1e>} imagemask} bind
{8 8 true tmpa {<df cf 8f 9f fd fc f8 f9>} imagemask} bind
{8 8 true tmpa {<ff 3f 3f ff ff f3 f3 ff>} imagemask} bind 7 array astore def
/ppaint { gsave clip tmpa dup setmatrix pathbbox neg exch neg 4 2 roll
  neg 4 -1 roll 2 copy gt {exch} if 8 div ceiling 8 mul 4 2 roll neg 2 copy
  gt {exch} if 8 div ceiling 8 mul 3 -1 roll -8 5 -1 roll
  { 3 index exch 5 exch put dup -8 3 index { 3 index
  exch 4 exch put 3 index exec } for } for pop pop pop pop grestore } bind def
/setstyles {
  currentlinewidth mul setlinewidth /style exch def
  style 1 and 0 gt not {closepath} if
  style 1024 and 0 gt {2 setlinecap} if
  style 2 and 0 gt {currentlinewidth 4 mul dup 2 array astore 0 setdash} if
  style 4 and 0 gt {0.5 currentlinewidth 4 mul 2 array astore 0 setdash} if
  gsave style 16 and 0 gt { style 224 and -5 bitshift style 256 and 0 gt {
  7 exch sub 8 div dup 1 exch sub currentrgbcolor 3 array astore
  {3 copy mul add 4 1 roll pop} forall pop pop setrgbcolor eofill}
  {dup 7 lt {gar exch get ppaint} {pop eofill} ifelse} ifelse}
  {style 256 and 0 gt {1 setgray eofill} if} ifelse grestore style 8 and 0 gt 
  style 512 eq or {newpath} {stroke} ifelse grestore} def     

/polygon { gsave /num exch def moveto num 1 sub {lineto} repeat setstyles } def
/xcarc   { gsave newpath arc setstyles } def
/elb { matrix currentmatrix 7 -1 roll 7 -1 roll translate 5 1 roll 4 -1 roll
	3 index div 1 scale } def
/ele { 0 4 1 roll 0 4 1 roll } bind def
/ellipse { gsave elb newpath ele arc setmatrix setstyles } def
/pellip  { elb ele arc setmatrix } def
/nellip  { elb ele arcn setmatrix } def
/spline  { gsave moveto curveto setstyles } def
/polyc   { {lineto} repeat } bind def
/beginpath { gsave moveto } bind def
/endpath { setstyles } bind def
/bop	 { 1 setlinecap 0 setlinejoin 6 setmiterlimit 0 0 0 scb cRedef } def
/psinsertion {/PSobj save def /showpage {} def /setpagedevice {pop} def bop
	rotate translate dup scale} def
/end_insert {PSobj restore} def
/setpagemat {/pagemat matrix currentmatrix def} def
/inchscale  {setpagemat 0.375 mul dup scale} def
/cmscale    {setpagemat 0.35433071 mul dup scale} def

%%EndResource
%%EndProlog

% XCircuit output starts here.

%%BeginSetup

/analog::source {
% hidden
begingate
1 1.000 0 0 32 0.000 360.000 xcarc
1 1.000 0 32 0 64 2 polygon
1 1.000 0 -32 0 -64 2 polygon
endgate
} def

/generic::arrowhead {
% nonetwork
begingate
8 -28 beginpath
3 -18 3 -15 0 0 curveto
-3 -15 -3 -18 -8 -28 curveto
-2 -26 2 -26 8 -28 curveto
249 
1.000 endpath
endgate
} def

/analog::isource {
begingate
1.000 0 0 0 analog::source
1 0.750 0 20 0 -8 2 polygon
0.800 180 0 -20 generic::arrowhead
1.000 0.000 0.000 scb
(i.p) {/Times-Roman cf} 2 9 0 1.000 0 64 pinlabel
(i.m) {/Times-Roman cf} 2 13 0 1.000 0 -64 pinlabel
endgate
} def

/analog::diode {
begingate
248 1.000 -18 -16 0 16 18 -16 3 polygon
1 1.000 0 -48 0 -16 2 polygon
1 1.000 0 48 0 16 2 polygon
1 1.000 -18 16 18 16 2 polygon
1.000 0.000 0.000 scb
(d.m) {/Times-Roman cf} 2 9 0 1.000 0 48 pinlabel
(d.p) {/Times-Roman cf} 2 13 0 1.000 0 -48 pinlabel
endgate
} def

/analog::gnd {
% trivial
begingate
1 1.000 0 0 0 -32 2 polygon
1 1.000 -32 -32 32 -32 2 polygon
1 1.000 -18 -46 18 -46 2 polygon
1 1.000 -4 -60 4 -60 2 polygon
0.933 0.604 0.000 scb
(GND) {/Times-Roman cf} 2 1 0 1.000 0 0 pinglobal
endgate
} def

/analog::vsource {
begingate
1.000 0 0 0 analog::source
(+) {/Symbol cf} 2 5 0 1.000 0 14 label
(-) {/Symbol cf} 2 5 0 1.000 0 -22 label
1.000 0.000 0.000 scb
(v.p) {/Times-Roman cf} 2 9 0 1.000 0 64 pinlabel
(v.m) {/Times-Roman cf} 2 13 0 1.000 0 -64 pinlabel
endgate
} def

/generic::dot {
% trivial
begingate
248 1.000 0 0 6 0.000 360.000 xcarc
1.000 0.000 0.000 scb
(x) {/Times-Roman cf} 2 29 0 1.000 0 0 pinlabel
endgate
} def


%%EndSetup

%%Page: XC4942.ttU1XB 1
%%PageOrientation: Portrait
/pgsave save def bop
1.0000 inchscale
2.6000 setlinewidth 960 476 translate

1.000 270 496 144 analog::isource
1.000 270 496 -96 analog::isource
1.000 270 -480 240 analog::isource
1.000 270 -480 0 analog::isource
1.000 270 -480 336 analog::diode
1.000 270 -480 80 analog::diode
1.000 270 496 224 analog::diode
1.000 270 496 -16 analog::diode
1.000 0 736 -224 analog::gnd
1.000 0 -416 -224 analog::gnd
1.000 90 -208 -32 analog::vsource
1.000 90 96 288 analog::vsource
1.000 90 -208 384 analog::vsource
1.000 90 -208 192 analog::vsource
1 1.000 -528 80 -528 0 -736 0 3 polygon
1 1.000 544 224 544 144 2 polygon
1 1.000 544 -16 544 -96 2 polygon
1.000 90 -96 384 analog::diode
1.000 90 -96 192 analog::diode
1.000 90 -96 -32 analog::diode
1 1.000 -416 240 -272 384 2 polygon
1 1.000 -416 240 -272 192 2 polygon
1 1.000 -416 240 -272 -32 2 polygon
1.000 90 96 96 analog::vsource
1.000 90 96 -128 analog::vsource
1 1.000 -416 0 -256 288 32 288 3 polygon
1 1.000 -416 0 -256 96 48 96 3 polygon
1.000 90 192 288 analog::diode
1.000 90 192 96 analog::diode
1.000 90 192 -128 analog::diode
1 1.000 240 -128 448 -96 2 polygon
1 1.000 -48 -32 240 -32 432 -96 3 polygon
1 1.000 -48 192 240 192 432 144 3 polygon
1 1.000 240 96 432 144 2 polygon
1 1.000 240 288 432 384 2 polygon
1 1.000 -48 384 432 384 2 polygon
1 1.000 560 144 736 144 2 polygon
1 1.000 560 -96 736 -96 2 polygon
1.000 0 -736 0 generic::dot
1.000 0 -416 0 generic::dot
1.000 0 -416 240 generic::dot
1.000 0 -528 240 generic::dot
1.000 0 -528 0 generic::dot
1.000 0 432 144 generic::dot
1.000 0 432 384 generic::dot
1.000 0 432 -96 generic::dot
1.000 0 544 -96 generic::dot
1.000 0 736 -96 generic::dot
1.000 0 736 144 generic::dot
1 1.000 448 224 432 224 432 144 3 polygon
1 1.000 448 -16 432 -16 432 -96 3 polygon
1 1.000 -416 240 -416 336 -432 336 3 polygon
1 1.000 -416 0 -416 80 -432 80 3 polygon
(v1) {/Helvetica cf} 2 16 0 1.000 208 208 label
(v2) {/Helvetica cf} 2 16 0 1.000 208 400 label
(v0) {/Helvetica cf} 2 16 0 1.000 208 -16 label
(7) {/Helvetica cf} 2 16 0 1.000 -224 432 label
(3) {/Helvetica cf} 2 16 0 1.000 -224 240 label
(2) {/Helvetica cf} 2 16 0 1.000 -224 16 label
(8) {/Helvetica cf} 2 16 0 1.000 80 336 label
(5) {/Helvetica cf} 2 16 0 1.000 80 144 label
(4) {/Helvetica cf} 2 16 0 1.000 80 -80 label
(1) {/Helvetica cf} 2 16 0 1.000 480 80 label
(1) {/Helvetica cf} 2 16 0 1.000 480 -160 label
(1) {/Helvetica cf} 2 16 0 1.000 -496 160 label
(1) {/Helvetica cf} 2 16 0 1.000 -496 -80 label
1 1.000 32 -128 -416 -128 2 polygon
1.000 180 -416 -176 analog::vsource
1.000 180 -272 -176 analog::vsource
1 1.000 -416 -112 -416 0 2 polygon
1 1.000 -272 -112 -272 -32 2 polygon
1.000 0 -272 -32 generic::dot
(u1) {/Helvetica cf} 2 16 0 1.000 -208 -176 label
(u0) {/Helvetica cf} 2 16 0 1.000 -512 -176 label
1.000 0 -272 -224 analog::gnd
1.000 0 -736 -224 analog::gnd
1 1.000 -528 336 -528 240 -736 240 -736 -240 4 polygon
0.000 0.000 0.000 scb
1.000 0 -416 -128 generic::dot
sce
1 1.000 432 384 736 384 736 -224 3 polygon
pgsave restore showpage

%%Trailer
XCIRCsave restore
%%EOF
